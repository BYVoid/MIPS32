library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Common.all;

entity Rom is
  port (
    addr: in Int10;
    data: out Int32
  );
end Rom;

architecture Behavioral of Rom is
  constant NUM_ROM_CELLS: integer := 1024;
  type RomType is array(0 to NUM_ROM_CELLS - 1) of Int32;
  signal rom: RomType;
begin
  data <= rom(to_integer(unsigned(addr)));
  rom(0) <= x"00000000";
  rom(1) <= x"10000001";
  rom(2) <= x"00000000";
  rom(3) <= x"3c08beff";
  rom(4) <= x"3508fff8";
  rom(5) <= x"240900ff";
  rom(6) <= x"ad090000";
  rom(7) <= x"3c10be00";
  rom(8) <= x"240f0000";
  rom(9) <= x"020f7821";
  rom(10) <= x"8de90000";
  rom(11) <= x"8def0004";
  rom(12) <= x"000f7c00";
  rom(13) <= x"012f4825";
  rom(14) <= x"3c08464c";
  rom(15) <= x"3508457f";
  rom(16) <= x"11090003";
  rom(17) <= x"00000000";
  rom(18) <= x"10000042";
  rom(19) <= x"00000000";
  rom(20) <= x"240f0038";
  rom(21) <= x"020f7821";
  rom(22) <= x"8df10000";
  rom(23) <= x"8def0004";
  rom(24) <= x"000f7c00";
  rom(25) <= x"022f8825";
  rom(26) <= x"240f0058";
  rom(27) <= x"020f7821";
  rom(28) <= x"8df20000";
  rom(29) <= x"8def0004";
  rom(30) <= x"000f7c00";
  rom(31) <= x"024f9025";
  rom(32) <= x"3252ffff";
  rom(33) <= x"240f0030";
  rom(34) <= x"020f7821";
  rom(35) <= x"8df30000";
  rom(36) <= x"8def0004";
  rom(37) <= x"000f7c00";
  rom(38) <= x"026f9825";
  rom(39) <= x"262f0008";
  rom(40) <= x"000f7840";
  rom(41) <= x"020f7821";
  rom(42) <= x"8df40000";
  rom(43) <= x"8def0004";
  rom(44) <= x"000f7c00";
  rom(45) <= x"028fa025";
  rom(46) <= x"262f0010";
  rom(47) <= x"000f7840";
  rom(48) <= x"020f7821";
  rom(49) <= x"8df50000";
  rom(50) <= x"8def0004";
  rom(51) <= x"000f7c00";
  rom(52) <= x"02afa825";
  rom(53) <= x"262f0004";
  rom(54) <= x"000f7840";
  rom(55) <= x"020f7821";
  rom(56) <= x"8df60000";
  rom(57) <= x"8def0004";
  rom(58) <= x"000f7c00";
  rom(59) <= x"02cfb025";
  rom(60) <= x"12800010";
  rom(61) <= x"00000000";
  rom(62) <= x"12a0000e";
  rom(63) <= x"00000000";
  rom(64) <= x"26cf0000";
  rom(65) <= x"000f7840";
  rom(66) <= x"020f7821";
  rom(67) <= x"8de80000";
  rom(68) <= x"8def0004";
  rom(69) <= x"000f7c00";
  rom(70) <= x"010f4025";
  rom(71) <= x"ae880000";
  rom(72) <= x"26d60004";
  rom(73) <= x"26940004";
  rom(74) <= x"26b5fffc";
  rom(75) <= x"1ea0fff4";
  rom(76) <= x"00000000";
  rom(77) <= x"26310020";
  rom(78) <= x"2652ffff";
  rom(79) <= x"1e40ffd7";
  rom(80) <= x"00000000";
  rom(81) <= x"02600008";
  rom(82) <= x"00000000";
  rom(83) <= x"1000ffff";
  rom(84) <= x"00000000";
  rom(85) <= x"1000ffff";
  rom(86) <= x"00000000";
end architecture;
