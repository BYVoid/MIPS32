library ieee;
use ieee.std_logic_1164.all;

entity CPU is
end CPU;

architecture Behavioral of CPU is

begin

end Behavioral;
